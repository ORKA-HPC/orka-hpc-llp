// Copyright (c) 2001-2018 Intel Corporation
//  
// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to
// permit persons to whom the Software is furnished to do so, subject to
// the following conditions:
//  
// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.
//  
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
// TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
// SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

`timescale 1 ps / 1 ps
`default_nettype none

// This is the top module of the design where the BSP is connected to external Pins
module a10_pcie_ref_design 
(
   //Dev Kit Pins
   output wire        board_pins_L0_led ,
   output wire        board_pins_alive_led , 
   output wire        board_pins_comp_led , 
   input wire         board_pins_free_clk , 
   output wire        board_pins_gen2_led , 
   output wire        board_pins_gen3_led , 
   output wire [ 3:0] board_pins_lane_active_led , 
   input wire         board_pins_req_compliance_pb , 
   input wire         board_pins_set_compliance_mode, 
   input wire         config_clk_clk , 
   input wire         pcie_rstn_npor , 
   input wire         pcie_rstn_pin_perst , 
   // DDR4
   input wire         pll_ref_clk , // reference clock for the DDR Memory PLL
   input wire         oct_rzqin ,
   output wire [ 1:0] mem_ba ,
   output wire [ 0:0] mem_bg ,
   output wire [ 0:0] mem_cke ,
   output wire [ 0:0] mem_ck ,
   output wire [ 0:0] mem_ck_n ,
   output wire [ 0:0] mem_cs_n ,
   output wire [ 0:0] mem_reset_n ,
   output wire [ 0:0] mem_odt ,
   output wire [ 0:0] mem_act_n ,
   output wire [16:0] mem_a ,
   inout wire [63:0]  mem_dq ,
   output wire [ 0:0] mem_par ,
   input wire [ 0:0]  mem_alert_n ,
   inout wire [ 7:0]  mem_dqs ,
   inout wire [ 7:0]  mem_dqs_n ,
   inout wire [ 7:0]  mem_dbi_n ,
   // PCIe
   input wire         ref_clk_clk , 
   input wire         xcvr_rx_in0 , 
   input wire         xcvr_rx_in1 , 
   input wire         xcvr_rx_in2 , 
   input wire         xcvr_rx_in3 , 
   input wire         xcvr_rx_in4 , 
   input wire         xcvr_rx_in5 , 
   input wire         xcvr_rx_in6 , 
   input wire         xcvr_rx_in7 , 
   output wire        xcvr_tx_out0 , 
   output wire        xcvr_tx_out1 , 
   output wire        xcvr_tx_out2 , 
   output wire        xcvr_tx_out3 , 
   output wire        xcvr_tx_out4 , 
   output wire        xcvr_tx_out5 , 
   output wire        xcvr_tx_out6 , 
   output wire        xcvr_tx_out7   
);
  

   bsp_top u_top 
   (
      // PLL 
      .pll_refclk_clk                                         ( config_clk_clk ),
      // DDR4 
      .ddr4_pll_ref_clk_clk                                   ( pll_ref_clk ),
      .ddr4_mem_mem_ck                                        ( mem_ck ),
      .ddr4_mem_mem_ck_n                                      ( mem_ck_n ),
      .ddr4_mem_mem_a                                         ( mem_a ),
      .ddr4_mem_mem_act_n                                     ( mem_act_n ),
      .ddr4_mem_mem_ba                                        ( mem_ba ),
      .ddr4_mem_mem_bg                                        ( mem_bg ),
      .ddr4_mem_mem_cke                                       ( mem_cke ),
      .ddr4_mem_mem_cs_n                                      ( mem_cs_n ),
      .ddr4_mem_mem_odt                                       ( mem_odt ),
      .ddr4_mem_mem_reset_n                                   ( mem_reset_n ),
      .ddr4_mem_mem_par                                       ( mem_par ),
      .ddr4_mem_mem_alert_n                                   ( mem_alert_n ),
      .ddr4_mem_mem_dqs                                       ( mem_dqs ),
      .ddr4_mem_mem_dqs_n                                     ( mem_dqs_n ),
      .ddr4_mem_mem_dq                                        ( mem_dq ),
      .ddr4_mem_mem_dbi_n                                     ( mem_dbi_n ),
      .ddr4_oct_oct_rzqin                                     ( oct_rzqin ),

      //Devkit
      .board_pins_L0_led                                      ( board_pins_L0_led ),
      .board_pins_alive_led                                   ( board_pins_alive_led ),
      .board_pins_comp_led                                    ( board_pins_comp_led ),
      .board_pins_free_clk                                    ( board_pins_free_clk ),
      .board_pins_gen2_led                                    ( board_pins_gen2_led ),
      .board_pins_gen3_led                                    ( board_pins_gen3_led ),
      .board_pins_lane_active_led                             ( board_pins_lane_active_led ),
      .board_pins_req_compliance_pb                           ( board_pins_req_compliance_pb ),
      .board_pins_set_compliance_mode                         ( board_pins_set_compliance_mode ),

      //PCIe 
      .a10_pcie_refclk_clk                                    ( ref_clk_clk ),
      .hip_ctrl_test_in                                       ( 0 ),
      .hip_ctrl_simu_mode_pipe                                ( 1'b0 ),
      .pcie_rstn_npor                                         ( pcie_rstn_npor ),
      .pcie_rstn_pin_perst                                    ( pcie_rstn_pin_perst ),
      .pipe_sim_only_sim_pipe_pclk_in                         ( 1'b0 ),
      .pipe_sim_only_sim_pipe_rate                            (),
      .pipe_sim_only_sim_ltssmstate                           (),
      .pipe_sim_only_eidleinfersel0                           (),
      .pipe_sim_only_eidleinfersel1                           (),
      .pipe_sim_only_eidleinfersel2                           (),
      .pipe_sim_only_eidleinfersel3                           (),
      .pipe_sim_only_eidleinfersel4                           (),
      .pipe_sim_only_eidleinfersel5                           (),
      .pipe_sim_only_eidleinfersel6                           (),
      .pipe_sim_only_eidleinfersel7                           (),
      .pipe_sim_only_powerdown0                               (),
      .pipe_sim_only_powerdown1                               (),
      .pipe_sim_only_powerdown2                               (),
      .pipe_sim_only_powerdown3                               (),
      .pipe_sim_only_powerdown4                               (),
      .pipe_sim_only_powerdown5                               (),
      .pipe_sim_only_powerdown6                               (),
      .pipe_sim_only_powerdown7                               (),
      .pipe_sim_only_rxpolarity0                              (),
      .pipe_sim_only_rxpolarity1                              (),
      .pipe_sim_only_rxpolarity2                              (),
      .pipe_sim_only_rxpolarity3                              (),
      .pipe_sim_only_rxpolarity4                              (),
      .pipe_sim_only_rxpolarity5                              (),
      .pipe_sim_only_rxpolarity6                              (),
      .pipe_sim_only_rxpolarity7                              (),
      .pipe_sim_only_txcompl0                                 (),
      .pipe_sim_only_txcompl1                                 (),
      .pipe_sim_only_txcompl2                                 (),
      .pipe_sim_only_txcompl3                                 (),
      .pipe_sim_only_txcompl4                                 (),
      .pipe_sim_only_txcompl5                                 (),
      .pipe_sim_only_txcompl6                                 (),
      .pipe_sim_only_txcompl7                                 (),
      .pipe_sim_only_txdata0                                  (),
      .pipe_sim_only_txdata1                                  (),
      .pipe_sim_only_txdata2                                  (),
      .pipe_sim_only_txdata3                                  (),
      .pipe_sim_only_txdata4                                  (),
      .pipe_sim_only_txdata5                                  (),
      .pipe_sim_only_txdata6                                  (),
      .pipe_sim_only_txdata7                                  (),
      .pipe_sim_only_txdatak0                                 (),
      .pipe_sim_only_txdatak1                                 (),
      .pipe_sim_only_txdatak2                                 (),
      .pipe_sim_only_txdatak3                                 (),
      .pipe_sim_only_txdatak4                                 (),
      .pipe_sim_only_txdatak5                                 (),
      .pipe_sim_only_txdatak6                                 (),
      .pipe_sim_only_txdatak7                                 (),
      .pipe_sim_only_txdetectrx0                              (),
      .pipe_sim_only_txdetectrx1                              (),
      .pipe_sim_only_txdetectrx2                              (),
      .pipe_sim_only_txdetectrx3                              (),
      .pipe_sim_only_txdetectrx4                              (),
      .pipe_sim_only_txdetectrx5                              (),
      .pipe_sim_only_txdetectrx6                              (),
      .pipe_sim_only_txdetectrx7                              (),
      .pipe_sim_only_txelecidle0                              (),
      .pipe_sim_only_txelecidle1                              (),
      .pipe_sim_only_txelecidle2                              (),
      .pipe_sim_only_txelecidle3                              (),
      .pipe_sim_only_txelecidle4                              (),
      .pipe_sim_only_txelecidle5                              (),
      .pipe_sim_only_txelecidle6                              (),
      .pipe_sim_only_txelecidle7                              (),
      .pipe_sim_only_txdeemph0                                (),
      .pipe_sim_only_txdeemph1                                (),
      .pipe_sim_only_txdeemph2                                (),
      .pipe_sim_only_txdeemph3                                (),
      .pipe_sim_only_txdeemph4                                (),
      .pipe_sim_only_txdeemph5                                (),
      .pipe_sim_only_txdeemph6                                (),
      .pipe_sim_only_txdeemph7                                (),
      .pipe_sim_only_txmargin0                                (),
      .pipe_sim_only_txmargin1                                (),
      .pipe_sim_only_txmargin2                                (),
      .pipe_sim_only_txmargin3                                (),
      .pipe_sim_only_txmargin4                                (),
      .pipe_sim_only_txmargin5                                (),
      .pipe_sim_only_txmargin6                                (),
      .pipe_sim_only_txmargin7                                (),
      .pipe_sim_only_txswing0                                 (),
      .pipe_sim_only_txswing1                                 (),
      .pipe_sim_only_txswing2                                 (),
      .pipe_sim_only_txswing3                                 (),
      .pipe_sim_only_txswing4                                 (),
      .pipe_sim_only_txswing5                                 (),
      .pipe_sim_only_txswing6                                 (),
      .pipe_sim_only_txswing7                                 (),
      .pipe_sim_only_phystatus0                               ( '0 ),
      .pipe_sim_only_phystatus1                               ( '0 ),
      .pipe_sim_only_phystatus2                               ( '0 ),
      .pipe_sim_only_phystatus3                               ( '0 ),
      .pipe_sim_only_phystatus4                               ( '0 ),
      .pipe_sim_only_phystatus5                               ( '0 ),
      .pipe_sim_only_phystatus6                               ( '0 ),
      .pipe_sim_only_phystatus7                               ( '0 ),
      .pipe_sim_only_rxdata0                                  ( '0 ),
      .pipe_sim_only_rxdata1                                  ( '0 ),
      .pipe_sim_only_rxdata2                                  ( '0 ),
      .pipe_sim_only_rxdata3                                  ( '0 ),
      .pipe_sim_only_rxdata4                                  ( '0 ),
      .pipe_sim_only_rxdata5                                  ( '0 ),
      .pipe_sim_only_rxdata6                                  ( '0 ),
      .pipe_sim_only_rxdata7                                  ( '0 ),
      .pipe_sim_only_rxdatak0                                 ( '0 ),
      .pipe_sim_only_rxdatak1                                 ( '0 ),
      .pipe_sim_only_rxdatak2                                 ( '0 ),
      .pipe_sim_only_rxdatak3                                 ( '0 ),
      .pipe_sim_only_rxdatak4                                 ( '0 ),
      .pipe_sim_only_rxdatak5                                 ( '0 ),
      .pipe_sim_only_rxdatak6                                 ( '0 ),
      .pipe_sim_only_rxdatak7                                 ( '0 ),
      .pipe_sim_only_rxelecidle0                              ( '0 ),
      .pipe_sim_only_rxelecidle1                              ( '0 ),
      .pipe_sim_only_rxelecidle2                              ( '0 ),
      .pipe_sim_only_rxelecidle3                              ( '0 ),
      .pipe_sim_only_rxelecidle4                              ( '0 ),
      .pipe_sim_only_rxelecidle5                              ( '0 ),
      .pipe_sim_only_rxelecidle6                              ( '0 ),
      .pipe_sim_only_rxelecidle7                              ( '0 ),
      .pipe_sim_only_rxstatus0                                ( '0 ),
      .pipe_sim_only_rxstatus1                                ( '0 ),
      .pipe_sim_only_rxstatus2                                ( '0 ),
      .pipe_sim_only_rxstatus3                                ( '0 ),
      .pipe_sim_only_rxstatus4                                ( '0 ),
      .pipe_sim_only_rxstatus5                                ( '0 ),
      .pipe_sim_only_rxstatus6                                ( '0 ),
      .pipe_sim_only_rxstatus7                                ( '0 ),
      .pipe_sim_only_rxvalid0                                 ( '0 ),
      .pipe_sim_only_rxvalid1                                 ( '0 ),
      .pipe_sim_only_rxvalid2                                 ( '0 ),
      .pipe_sim_only_rxvalid3                                 ( '0 ),
      .pipe_sim_only_rxvalid4                                 ( '0 ),
      .pipe_sim_only_rxvalid5                                 ( '0 ),
      .pipe_sim_only_rxvalid6                                 ( '0 ),
      .pipe_sim_only_rxvalid7                                 ( '0 ),
      .pipe_sim_only_rxdataskip0                              ( '0 ),
      .pipe_sim_only_rxdataskip1                              ( '0 ),
      .pipe_sim_only_rxdataskip2                              ( '0 ),
      .pipe_sim_only_rxdataskip3                              ( '0 ),
      .pipe_sim_only_rxdataskip4                              ( '0 ),
      .pipe_sim_only_rxdataskip5                              ( '0 ),
      .pipe_sim_only_rxdataskip6                              ( '0 ),
      .pipe_sim_only_rxdataskip7                              ( '0 ),
      .pipe_sim_only_rxblkst0                                 ( '0 ),
      .pipe_sim_only_rxblkst1                                 ( '0 ),
      .pipe_sim_only_rxblkst2                                 ( '0 ),
      .pipe_sim_only_rxblkst3                                 ( '0 ),
      .pipe_sim_only_rxblkst4                                 ( '0 ),
      .pipe_sim_only_rxblkst5                                 ( '0 ),
      .pipe_sim_only_rxblkst6                                 ( '0 ),
      .pipe_sim_only_rxblkst7                                 ( '0 ),
      .pipe_sim_only_rxsynchd0                                ( '0 ),
      .pipe_sim_only_rxsynchd1                                ( '0 ),
      .pipe_sim_only_rxsynchd2                                ( '0 ),
      .pipe_sim_only_rxsynchd3                                ( '0 ),
      .pipe_sim_only_rxsynchd4                                ( '0 ),
      .pipe_sim_only_rxsynchd5                                ( '0 ),
      .pipe_sim_only_rxsynchd6                                ( '0 ),
      .pipe_sim_only_rxsynchd7                                ( '0 ),
      .pipe_sim_only_currentcoeff0                            (),
      .pipe_sim_only_currentcoeff1                            (),
      .pipe_sim_only_currentcoeff2                            (),
      .pipe_sim_only_currentcoeff3                            (),
      .pipe_sim_only_currentcoeff4                            (),
      .pipe_sim_only_currentcoeff5                            (),
      .pipe_sim_only_currentcoeff6                            (),
      .pipe_sim_only_currentcoeff7                            (),
      .pipe_sim_only_currentrxpreset0                         (),
      .pipe_sim_only_currentrxpreset1                         (),
      .pipe_sim_only_currentrxpreset2                         (),
      .pipe_sim_only_currentrxpreset3                         (),
      .pipe_sim_only_currentrxpreset4                         (),
      .pipe_sim_only_currentrxpreset5                         (),
      .pipe_sim_only_currentrxpreset6                         (),
      .pipe_sim_only_currentrxpreset7                         (),
      .pipe_sim_only_txsynchd0                                (),
      .pipe_sim_only_txsynchd1                                (),
      .pipe_sim_only_txsynchd2                                (),
      .pipe_sim_only_txsynchd3                                (),
      .pipe_sim_only_txsynchd4                                (),
      .pipe_sim_only_txsynchd5                                (),
      .pipe_sim_only_txsynchd6                                (),
      .pipe_sim_only_txsynchd7                                (),
      .pipe_sim_only_txblkst0                                 (),
      .pipe_sim_only_txblkst1                                 (),
      .pipe_sim_only_txblkst2                                 (),
      .pipe_sim_only_txblkst3                                 (),
      .pipe_sim_only_txblkst4                                 (),
      .pipe_sim_only_txblkst5                                 (),
      .pipe_sim_only_txblkst6                                 (),
      .pipe_sim_only_txblkst7                                 (),
      .pipe_sim_only_txdataskip0                              (),
      .pipe_sim_only_txdataskip1                              (),
      .pipe_sim_only_txdataskip2                              (),
      .pipe_sim_only_txdataskip3                              (),
      .pipe_sim_only_txdataskip4                              (),
      .pipe_sim_only_txdataskip5                              (),
      .pipe_sim_only_txdataskip6                              (),
      .pipe_sim_only_txdataskip7                              (),
      .pipe_sim_only_rate0                                    (),
      .pipe_sim_only_rate1                                    (),
      .pipe_sim_only_rate2                                    (),
      .pipe_sim_only_rate3                                    (),
      .pipe_sim_only_rate4                                    (),
      .pipe_sim_only_rate5                                    (),
      .pipe_sim_only_rate6                                    (),
      .pipe_sim_only_rate7                                    (),
      .xcvr_rx_in0                                            ( xcvr_rx_in0 ),
      .xcvr_rx_in1                                            ( xcvr_rx_in1 ),
      .xcvr_rx_in2                                            ( xcvr_rx_in2 ),
      .xcvr_rx_in3                                            ( xcvr_rx_in3 ),
      .xcvr_rx_in4                                            ( xcvr_rx_in4 ),
      .xcvr_rx_in5                                            ( xcvr_rx_in5 ),
      .xcvr_rx_in6                                            ( xcvr_rx_in6 ),
      .xcvr_rx_in7                                            ( xcvr_rx_in7 ),
      .xcvr_tx_out0                                           ( xcvr_tx_out0 ),
      .xcvr_tx_out1                                           ( xcvr_tx_out1 ),
      .xcvr_tx_out2                                           ( xcvr_tx_out2 ),
      .xcvr_tx_out3                                           ( xcvr_tx_out3 ),
      .xcvr_tx_out4                                           ( xcvr_tx_out4 ),
      .xcvr_tx_out5                                           ( xcvr_tx_out5 ),
      .xcvr_tx_out6                                           ( xcvr_tx_out6 ),
      .xcvr_tx_out7                                           ( xcvr_tx_out7 )
   );

   

endmodule
